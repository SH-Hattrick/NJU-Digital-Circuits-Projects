module RAM2(
);


endmodule 